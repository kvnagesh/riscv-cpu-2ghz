//==============================================================================
// Copyright (c) 2025 Nagesh Vishnumurthy
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//==============================================================================

//==============================================================================
// File: riscv_ex3_stage.sv
// Description: Execute Stage 3 (EX3) - Stage 5 of 10 - RV64I Support
// Purpose: ALU computation stage 2, data forwarding (64-bit)
// Critical Path: < 500ps for 2 GHz @ 7nm
//==============================================================================

module riscv_ex3_stage (
    input  logic        clk,
    input  logic        rst_n,
    
    // Inputs from EX2 Stage
    input  logic [63:0] ex2_pc,
    input  logic [31:0] ex2_inst,
    input  logic [63:0] ex2_alu_result,
    input  logic [63:0] ex2_rs2_data,
    input  logic [4:0]  ex2_rd_addr,
    input  logic [2:0]  ex2_funct3,
    input  logic        ex2_valid,
    
    // Outputs to EX4 Stage - Pipeline Registers
    output logic [63:0] ex3_pc,         // NO RESET - Data path
    output logic [31:0] ex3_inst,       // NO RESET - Data path
    output logic [63:0] ex3_alu_result, // NO RESET - Data path (64-bit)
    output logic [63:0] ex3_rs2_data,   // NO RESET - Data path (64-bit)
    output logic [4:0]  ex3_rd_addr,    // NO RESET - Data path
    output logic [2:0]  ex3_funct3,     // NO RESET - Data path
    output logic        ex3_valid       // WITH RESET - Control path
);

    //==========================================================================
    // Pipeline Registers - NO RESET (Data Path)
    //==========================================================================
    always_ff @(posedge clk) begin
        ex3_pc         <= ex2_pc;
        ex3_inst       <= ex2_inst;
        ex3_alu_result <= ex2_alu_result;
        ex3_rs2_data   <= ex2_rs2_data;
        ex3_rd_addr    <= ex2_rd_addr;
        ex3_funct3     <= ex2_funct3;
    end
    
    //==========================================================================
    // Valid Signal - WITH RESET (Control Path)
    //==========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            ex3_valid <= 1'b0;
        else
            ex3_valid <= ex2_valid;
    end

endmodule
